
`define DATA_WIDTH 64 

`define PIXEL_IN_WIDTH 8 
`define PIXEL_OUT_WIDTH 8 

`define NUM_PIXEL_CHANEL_IN 8
`define NUM_PIXEL_CHANEL_OUT 8

`define WIDTH_FRAME 640 
`define HEIGHT_FRAME 480 

`define WIDTH_FIFO `DATA_WIDTH
`define NUM_WORDS_FIFO `WIDTH_FRAME*`HEIGHT_FRAME*`PIXEL_IN_WIDTH/`DATA_WIDTH
`define LOG2_NUM_WORDS_FIFO $clog2(`NUM_WORDS_FIFO)

`define NUM_WORDS_LINE_DILATE `WIDTH_FRAME / `NUM_PIXEL_CHANEL_IN

`define NUM_WORDS_CHANEL_IN  `NUM_WORDS_FIFO
`define NUM_WORDS_CHANEL_OUT `NUM_WORDS_FIFO

`define RANGE_DIFFERENCE 2